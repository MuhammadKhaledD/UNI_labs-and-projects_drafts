module seven_seg (I, S);

    input [11:0] I;
    output reg [20:0] S;

    reg [3:0] i [2:0];
    reg [6:0] s [2:0];
    integer j;

    always @(*) begin
        s[0] = 7'b1111111;
        s[1] = 7'b1111111;
        s[2] = 7'b1111111;

        i[2] = I[11:8];
        i[1] = I[7:4];
        i[0] = I[3:0];

        for (j = 2; j >= 0; j = j - 1) begin
            s[j][0] = (i[j][0] & ~i[j][1] & ~i[j][2] & ~i[j][3] | ~i[j][0] & ~i[j][1] & i[j][2] & ~i[j][3]);
            s[j][1] = (i[j][0] & ~i[j][1] & i[j][2] & ~i[j][3] | ~i[j][0] & i[j][1] & i[j][2] & ~i[j][3]);
            s[j][2] = ~i[j][0] & i[j][1] & ~i[j][2] & ~i[j][3];
            s[j][3] = (i[j][2] & i[j][0] & i[j][1] | i[j][2] & ~i[j][0] & ~i[j][1] | i[j][0] & ~i[j][1] & ~i[j][2] & ~i[j][3]);
            s[j][4] = (i[j][0] | ~i[j][1] & i[j][2]);
            s[j][5] = (i[j][0] & i[j][1] | i[j][1] & ~i[j][2] & ~i[j][3] | i[j][0] & ~i[j][2] & ~i[j][3]);
            s[j][6] = (~i[j][1] & ~i[j][2] & ~i[j][3] | i[j][0] & i[j][1] & i[j][2]);
        end

        S = {s[2], s[1], s[0]};
    end

endmodule