module display_controller(
    input [8:0] value,
    output [6:0] hex0,
    output [6:0] hex1,
    output [6:0] hex2
);
    wire [3:0] bcd0, bcd1, bcd2;
    
    // Convert binary to BCD
    binary_to_bcd bcd_converter(
        .binary(value),
        .bcd0(bcd0),
        .bcd1(bcd1),
        .bcd2(bcd2)
    );
    
    // Convert BCD to seven segment
    seven_segment_decoder seg0(
        .bin(bcd0),
        .seg(hex0)
    );
    
    seven_segment_decoder seg1(
        .bin(bcd1),
        .seg(hex1)
    );
    
    seven_segment_decoder seg2(
        .bin(bcd2),
        .seg(hex2)
    );
endmodule